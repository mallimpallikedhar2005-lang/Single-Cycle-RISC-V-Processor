module program_counter(clk,reset,pc_next,pc);
input clk, reset;
input [31:0] pc_next;
output reg [31:0] pc;
always @ (posedge clk or posedge reset)
begin
if (reset)
     pc <= 32'b0;
else 
  pc <= pc_next;
end
endmodule 