module AND_gate(input Branch,
                  input zero,
                  output out );
assign out = Branch & zero;
endmodule
